class fifo_env extends uvm_env;

endclass : fifo_env
