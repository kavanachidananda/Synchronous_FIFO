class fifo-seq_item extends uvm_sequence_item;
