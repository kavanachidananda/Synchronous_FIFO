class fifo_passive_agent extends uvm_agent;

endclass : fifo_passive_agent
