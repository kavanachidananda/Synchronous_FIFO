class fifo_scoreboard extends uvm_scoreboard;

endclass : fifo_scoreboard
