class fifo_sequence extends sequence #(fifo_transaction)
