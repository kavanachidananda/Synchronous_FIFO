`include "fifo_output_monitor.sv"

class fifo_passive_agent extends uvm_agent;
  fifo_output_monitor o_mon;
  'uvm_component_utils("fifo_passive_agent")

  function
endclass : fifo_passive_agent
