class fifo_test extends uvm_test;
endclass : fifo_test
