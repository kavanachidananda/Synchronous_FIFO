class fifo_driver extends uvm_driver #(fifo_sequence_item);

endclass : fifo_driver
